//
// Template for UVM-compliant configuration class
//

`ifndef RVV_FIFO_CFG__SV
`define RVV_FIFO_CFG__SV

class rvv_fifo_cfg extends uvm_object; 

   // Define test configuration parameters (e.g. how long to run)
   rand int num_trans;
   rand int num_scen;
   // ToDo: Add other environment configuration varaibles

   constraint cst_num_trans_default {
      num_trans inside {[1:7]};
   }
   constraint cst_num_scen_default {
      num_scen inside {[1:2]};
   }
   // ToDo: Add constraint blocks to prevent error injection

   `uvm_object_utils_begin(rvv_fifo_cfg)
      `uvm_field_int(num_trans,UVM_ALL_ON) 
      `uvm_field_int(num_scen,UVM_ALL_ON)
      // ToDo: add properties using macros here

   `uvm_object_utils_end

   extern function new(string name = "");
  
endclass: rvv_fifo_cfg

function rvv_fifo_cfg::new(string name = "");
   super.new(name);
endfunction: new


`endif // RVV_FIFO_CFG__SV
