
typedef enum logic [0:0]{
  ADDSUB_VADD, 
  ADDSUB_VSUB
} F_ADDSUB_t;               
