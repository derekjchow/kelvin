`ifndef RVV_CONFIG_SVH
`define RVV_CONFIG_SVH

`define ASSERT_ON

`endif // RVV_CONFIG_SVH