`ifndef RVV_CONFIG_SVH
`define RVV_CONFIG_SVH


//`define MULTI_LSU
`define MULTI_ALU
`define MULTI_MUL
`define MULTI_PMTRDT
//`define MULTI_DIV

`endif // RVV_CONFIG_SVH