// 31 down to 0
128'hffff0001ffff0002ffff0003ffff001f,
128'hffff0001ffff0002ffff0003ffff001e,
128'hffff0001ffff0002ffff0003ffff001d,
128'hffff0001ffff0002ffff0003ffff001c,
128'hffff0001ffff0002ffff0003ffff001b,
128'hffff0001ffff0002ffff0003ffff001a,
128'hffff0001ffff0002ffff0003ffff0019,
128'hffff0001ffff0002ffff0003ffff0018,
128'hffff0001ffff0002ffff0003ffff0017,
128'hffff0001ffff0002ffff0003ffff0016,
128'hffff0001ffff0002ffff0003ffff0015,
128'hffff0001ffff0002ffff0003ffff0014,
128'hffff0001ffff0002ffff0003ffff0013,
128'hffff0001ffff0002ffff0003ffff0012,
128'hffff0001ffff0002ffff0003ffff0011,
128'hffff0001ffff0002ffff0003ffff0010,
128'hffff0001ffff0002ffff0003ffff000f,
128'hffff0001ffff0002ffff0003ffff000e,
128'hffff0001ffff0002ffff0003ffff000d,
128'hffff0001ffff0002ffff0003ffff000c,
128'hffff0001ffff0002ffff0003ffff000b,
128'hffff0001ffff0002ffff0003ffff000a,
128'hffff0001ffff0002ffff0003ffff0009,
128'hffff0001ffff0002ffff0003ffff0008,
128'hffff0001ffff0002ffff0003ffff0007,
128'hffff0001ffff0002ffff0003ffff0006,
128'hffff0001ffff0002ffff0003ffff0005,
128'hffff0001ffff0002ffff0003ffff0004,
128'hffff0001ffff0002ffff0003ffff0003,
128'hffff0001ffff0002ffff0003ffff0001,
128'h0
