`ifndef RVV_CONFIG_SVH
`define RVV_CONFIG_SVH

// config for multi-issue
`define ISSUE_3_READ_PORT_6
//`define ISSUE_2_READ_PORT_6
//`define ISSUE_2_READ_PORT_4

`endif // RVV_CONFIG_SVH
