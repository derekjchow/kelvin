typedef enum logic [0:0]{
  ADDSUB_VADD, 
  ADDSUB_VSUB
} F_ADDSUB_t;   

typedef enum logic [1:0]{
  SHIFT_SLL, 
  SHIFT_SRL,
  SHIFT_SRA
} F_SHIFT_t;   

