`ifndef RVV_BACKEND_TB_SV
`define RVV_BACKEND_TB_SV

`include "mstr_slv_src.incl"
`include "mstr_slv_intfs.incl"

`include "rvv_cfg.sv"


`include "rvv_scoreboard.sv"

`include "rvv_cov.sv"

`endif // RVV_BACKEND_TB__SV
