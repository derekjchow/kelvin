// Copyright 2025 Google LLC
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.

//----------------------------------------------------------------------------
// Description:covergroup for RV32I instruction
//----------------------------------------------------------------------------
covergroup cvgrp_RV32_I;

	option.per_instance = 1;

	// base cover
	add: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {ADD};
		option.weight = 1;
	 }

	sub: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {SUB};
		option.weight = 1;
	 }

	cp_xor: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {XOR};
		option.weight = 1;
	 }

	cp_or: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {OR};
		option.weight = 1;
	 }

	cp_and: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {AND};
		option.weight = 1;
	 }

	sll: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {SLL};
		option.weight = 1;
	 }

	srl: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {SRL};
		option.weight = 1;
	 }

	sra: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {SRA};
		option.weight = 1;
	 }

	slt: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {SLT};
		option.weight = 1;
	 }

	sltu: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {SLTU};
		option.weight = 1;
	 }

	addi: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {ADDI};
		option.weight = 1;
	 }

	xori: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {XORI};
		option.weight = 1;
	 }

	ori: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {ORI};
		option.weight = 1;
	 }

	andi: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {ANDI};
		option.weight = 1;
	 }

	slli: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {SLLI};
		option.weight = 1;
	 }

	srli: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {SRLI};
		option.weight = 1;
	 }

	srai: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {SRAI};
		option.weight = 1;
	 }

	slti: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {SLTI};
		option.weight = 1;
	 }

	sltiu: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {SLTIU};
		option.weight = 1;
	 }

	lb: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {LB};
		option.weight = 1;
	 }

	lh: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {LH};
		option.weight = 1;
	 }

	lw: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {LW};
		option.weight = 1;
	 }

	lbu: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {LBU};
		option.weight = 1;
	 }

	lhu: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {LHU};
		option.weight = 1;
	 }

	sb: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {SB};
		option.weight = 1;
	 }

	sh: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {SH};
		option.weight = 1;
	 }

	sw: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {SW};
		option.weight = 1;
	 }

	beq: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {BEQ};
		option.weight = 1;
	 }

	bne: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {BNE};
		option.weight = 1;
	 }

	blt: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {BLT};
		option.weight = 1;
	 }

	bge: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {BGE};
		option.weight = 1;
	 }

	bltu: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {BLTU};
		option.weight = 1;
	 }

	bgeu: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {BGEU};
		option.weight = 1;
	 }

	jal: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {JAL};
		option.weight = 1;
	 }

	jalr: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {JALR};
		option.weight = 1;
	 }

	lui: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {LUI};
		option.weight = 1;
	 }

	auipc: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {AUIPC};
		option.weight = 1;
	 }

	ecall: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {ECALL};
		option.weight = 1;
	 }

	ebreak: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {EBREAK};
		option.weight = 1;
	 }

	fence: coverpoint rv32i_trans.insn_name iff(rv32i_trans.trap==0) {
		bins b0 = {FENCE};
		option.weight = 1;
	 }

	//RD (GPR) register assignment,x0 always 0
	rd_addr: coverpoint rv32i_trans.rd_addr iff(rv32i_trans.trap==0) {
		bins b0 = {0};
		bins b1 = {1};
		bins b2 = {2};
		bins b3 = {3};
		bins b4 = {4};
		bins b5 = {5};
		bins b6 = {6};
		bins b7 = {7};
		bins b8 = {8};
		bins b9 = {9};
		bins b10 = {10};
		bins b11 = {11};
		bins b12 = {12};
		bins b13 = {13};
		bins b14 = {14};
		bins b15 = {15};
		bins b16 = {16};
		bins b17 = {17};
		bins b18 = {18};
		bins b19 = {19};
		bins b20 = {20};
		bins b21 = {21};
		bins b22 = {22};
		bins b23 = {23};
		bins b24 = {24};
		bins b25 = {25};
		bins b26 = {26};
		bins b27 = {27};
		bins b28 = {28};
		bins b29 = {29};
		bins b30 = {30};
		bins b31 = {31};
		option.weight = 1;
	 }

	//RS1 (GPR) register assignment
	rs1_addr: coverpoint rv32i_trans.rs1_addr iff(rv32i_trans.trap==0) {
		bins b0 = {0};
		bins b1 = {1};
		bins b2 = {2};
		bins b3 = {3};
		bins b4 = {4};
		bins b5 = {5};
		bins b6 = {6};
		bins b7 = {7};
		bins b8 = {8};
		bins b9 = {9};
		bins b10 = {10};
		bins b11 = {11};
		bins b12 = {12};
		bins b13 = {13};
		bins b14 = {14};
		bins b15 = {15};
		bins b16 = {16};
		bins b17 = {17};
		bins b18 = {18};
		bins b19 = {19};
		bins b20 = {20};
		bins b21 = {21};
		bins b22 = {22};
		bins b23 = {23};
		bins b24 = {24};
		bins b25 = {25};
		bins b26 = {26};
		bins b27 = {27};
		bins b28 = {28};
		bins b29 = {29};
		bins b30 = {30};
		bins b31 = {31};
		option.weight = 1;
	 }

	//RS2 (GPR) register assignment
	rs2_addr: coverpoint rv32i_trans.rs2_addr iff(rv32i_trans.trap==0) {
		bins b0 = {0};
		bins b1 = {1};
		bins b2 = {2};
		bins b3 = {3};
		bins b4 = {4};
		bins b5 = {5};
		bins b6 = {6};
		bins b7 = {7};
		bins b8 = {8};
		bins b9 = {9};
		bins b10 = {10};
		bins b11 = {11};
		bins b12 = {12};
		bins b13 = {13};
		bins b14 = {14};
		bins b15 = {15};
		bins b16 = {16};
		bins b17 = {17};
		bins b18 = {18};
		bins b19 = {19};
		bins b20 = {20};
		bins b21 = {21};
		bins b22 = {22};
		bins b23 = {23};
		bins b24 = {24};
		bins b25 = {25};
		bins b26 = {26};
		bins b27 = {27};
		bins b28 = {28};
		bins b29 = {29};
		bins b30 = {30};
		bins b31 = {31};
		option.weight = 1;
	 }

	//RD toggle bits
	rd_val: coverpoint unsigned'(rv32i_trans.rd_val) iff(rv32i_trans.trap==0) {
		wildcard bins b_1_0_0 	= (32'b???????????????????????????????1=>32'b???????????????????????????????0);
		wildcard bins b_1_0_1 	= (32'b??????????????????????????????1?=>32'b??????????????????????????????0?);
		wildcard bins b_1_0_2 	= (32'b?????????????????????????????1??=>32'b?????????????????????????????0??);
		wildcard bins b_1_0_3 	= (32'b????????????????????????????1???=>32'b????????????????????????????0???);
		wildcard bins b_1_0_4 	= (32'b???????????????????????????1????=>32'b???????????????????????????0????);
		wildcard bins b_1_0_5 	= (32'b??????????????????????????1?????=>32'b??????????????????????????0?????);
		wildcard bins b_1_0_6 	= (32'b?????????????????????????1??????=>32'b?????????????????????????0??????);
		wildcard bins b_1_0_7 	= (32'b????????????????????????1???????=>32'b????????????????????????0???????);
		wildcard bins b_1_0_8 	= (32'b???????????????????????1????????=>32'b???????????????????????0????????);
		wildcard bins b_1_0_9 	= (32'b??????????????????????1?????????=>32'b??????????????????????0?????????);
		wildcard bins b_1_0_10 	= (32'b?????????????????????1??????????=>32'b?????????????????????0??????????);
		wildcard bins b_1_0_11 	= (32'b????????????????????1???????????=>32'b????????????????????0???????????);
		wildcard bins b_1_0_12 	= (32'b???????????????????1????????????=>32'b???????????????????0????????????);
		wildcard bins b_1_0_13 	= (32'b??????????????????1?????????????=>32'b??????????????????0?????????????);
		wildcard bins b_1_0_14 	= (32'b?????????????????1??????????????=>32'b?????????????????0??????????????);
		wildcard bins b_1_0_15 	= (32'b????????????????1???????????????=>32'b????????????????0???????????????);
		wildcard bins b_1_0_16 	= (32'b???????????????1????????????????=>32'b???????????????0????????????????);
		wildcard bins b_1_0_17 	= (32'b??????????????1?????????????????=>32'b??????????????0?????????????????);
		wildcard bins b_1_0_18 	= (32'b?????????????1??????????????????=>32'b?????????????0??????????????????);
		wildcard bins b_1_0_19 	= (32'b????????????1???????????????????=>32'b????????????0???????????????????);
		wildcard bins b_1_0_20 	= (32'b???????????1????????????????????=>32'b???????????0????????????????????);
		wildcard bins b_1_0_21 	= (32'b??????????1?????????????????????=>32'b??????????0?????????????????????);
		wildcard bins b_1_0_22 	= (32'b?????????1??????????????????????=>32'b?????????0??????????????????????);
		wildcard bins b_1_0_23 	= (32'b????????1???????????????????????=>32'b????????0???????????????????????);
		wildcard bins b_1_0_24 	= (32'b???????1????????????????????????=>32'b???????0????????????????????????);
		wildcard bins b_1_0_25 	= (32'b??????1?????????????????????????=>32'b??????0?????????????????????????);
		wildcard bins b_1_0_26 	= (32'b?????1??????????????????????????=>32'b?????0??????????????????????????);
		wildcard bins b_1_0_27 	= (32'b????1???????????????????????????=>32'b????0???????????????????????????);
		wildcard bins b_1_0_28 	= (32'b???1????????????????????????????=>32'b???0????????????????????????????);
		wildcard bins b_1_0_29 	= (32'b??1?????????????????????????????=>32'b??0?????????????????????????????);
		wildcard bins b_1_0_30 	= (32'b?1??????????????????????????????=>32'b?0??????????????????????????????);
		wildcard bins b_1_0_31 	= (32'b1???????????????????????????????=>32'b0???????????????????????????????);
		wildcard bins b_0_1_0 	= (32'b???????????????????????????????0=>32'b???????????????????????????????1);
		wildcard bins b_0_1_1 	= (32'b??????????????????????????????0?=>32'b??????????????????????????????1?);
		wildcard bins b_0_1_2 	= (32'b?????????????????????????????0??=>32'b?????????????????????????????1??);
		wildcard bins b_0_1_3 	= (32'b????????????????????????????0???=>32'b????????????????????????????1???);
		wildcard bins b_0_1_4 	= (32'b???????????????????????????0????=>32'b???????????????????????????1????);
		wildcard bins b_0_1_5 	= (32'b??????????????????????????0?????=>32'b??????????????????????????1?????);
		wildcard bins b_0_1_6 	= (32'b?????????????????????????0??????=>32'b?????????????????????????1??????);
		wildcard bins b_0_1_7 	= (32'b????????????????????????0???????=>32'b????????????????????????1???????);
		wildcard bins b_0_1_8 	= (32'b???????????????????????0????????=>32'b???????????????????????1????????);
		wildcard bins b_0_1_9 	= (32'b??????????????????????0?????????=>32'b??????????????????????1?????????);
		wildcard bins b_0_1_10 	= (32'b?????????????????????0??????????=>32'b?????????????????????1??????????);
		wildcard bins b_0_1_11 	= (32'b????????????????????0???????????=>32'b????????????????????1???????????);
		wildcard bins b_0_1_12 	= (32'b???????????????????0????????????=>32'b???????????????????1????????????);
		wildcard bins b_0_1_13 	= (32'b??????????????????0?????????????=>32'b??????????????????1?????????????);
		wildcard bins b_0_1_14 	= (32'b?????????????????0??????????????=>32'b?????????????????1??????????????);
		wildcard bins b_0_1_15 	= (32'b????????????????0???????????????=>32'b????????????????1???????????????);
		wildcard bins b_0_1_16 	= (32'b???????????????0????????????????=>32'b???????????????1????????????????);
		wildcard bins b_0_1_17 	= (32'b??????????????0?????????????????=>32'b??????????????1?????????????????);
		wildcard bins b_0_1_18 	= (32'b?????????????0??????????????????=>32'b?????????????1??????????????????);
		wildcard bins b_0_1_19 	= (32'b????????????0???????????????????=>32'b????????????1???????????????????);
		wildcard bins b_0_1_20 	= (32'b???????????0????????????????????=>32'b???????????1????????????????????);
		wildcard bins b_0_1_21 	= (32'b??????????0?????????????????????=>32'b??????????1?????????????????????);
		wildcard bins b_0_1_22 	= (32'b?????????0??????????????????????=>32'b?????????1??????????????????????);
		wildcard bins b_0_1_23 	= (32'b????????0???????????????????????=>32'b????????1???????????????????????);
		wildcard bins b_0_1_24 	= (32'b???????0????????????????????????=>32'b???????1????????????????????????);
		wildcard bins b_0_1_25 	= (32'b??????0?????????????????????????=>32'b??????1?????????????????????????);
		wildcard bins b_0_1_26 	= (32'b?????0??????????????????????????=>32'b?????1??????????????????????????);
		wildcard bins b_0_1_27 	= (32'b????0???????????????????????????=>32'b????1???????????????????????????);
		wildcard bins b_0_1_28 	= (32'b???0????????????????????????????=>32'b???1????????????????????????????);
		wildcard bins b_0_1_29 	= (32'b??0?????????????????????????????=>32'b??1?????????????????????????????);
		wildcard bins b_0_1_30 	= (32'b?0??????????????????????????????=>32'b?1??????????????????????????????);
		wildcard bins b_0_1_31 	= (32'b0???????????????????????????????=>32'b1???????????????????????????????);
		option.weight = 1;
	 }

	//RD special values
	rd_sp_val: coverpoint unsigned'(rv32i_trans.rd_val) iff(rv32i_trans.trap==0) {
		bins b0 = {32'b0};
		bins b1 = {32'b00000000000000000000000000000001};
		bins b2 = {32'b11111111111111111111111111111111};
		bins b3 = {32'b01111111111111111111111111111111};
		bins b4 = {32'b10000000000000000000000000000000};
		bins b5 = {32'b10000000000000000000000000000001};
		option.weight = 1;
	 }

	//RD value sign
	rd_val_sign: coverpoint rv32i_trans.rd_val iff(rv32i_trans.trap==0) {
		bins b0 = {[$:-1]};
		bins b1 = {[1:$]};
		option.weight = 1;
	 }

	//RS1 toggle bits
	rs1_val: coverpoint unsigned'(rv32i_trans.rs1_val) iff(rv32i_trans.trap==0) {
		wildcard bins b_1_0_0 	= (32'b???????????????????????????????1=>32'b???????????????????????????????0);
		wildcard bins b_1_0_1 	= (32'b??????????????????????????????1?=>32'b??????????????????????????????0?);
		wildcard bins b_1_0_2 	= (32'b?????????????????????????????1??=>32'b?????????????????????????????0??);
		wildcard bins b_1_0_3 	= (32'b????????????????????????????1???=>32'b????????????????????????????0???);
		wildcard bins b_1_0_4 	= (32'b???????????????????????????1????=>32'b???????????????????????????0????);
		wildcard bins b_1_0_5 	= (32'b??????????????????????????1?????=>32'b??????????????????????????0?????);
		wildcard bins b_1_0_6 	= (32'b?????????????????????????1??????=>32'b?????????????????????????0??????);
		wildcard bins b_1_0_7 	= (32'b????????????????????????1???????=>32'b????????????????????????0???????);
		wildcard bins b_1_0_8 	= (32'b???????????????????????1????????=>32'b???????????????????????0????????);
		wildcard bins b_1_0_9 	= (32'b??????????????????????1?????????=>32'b??????????????????????0?????????);
		wildcard bins b_1_0_10 	= (32'b?????????????????????1??????????=>32'b?????????????????????0??????????);
		wildcard bins b_1_0_11 	= (32'b????????????????????1???????????=>32'b????????????????????0???????????);
		wildcard bins b_1_0_12 	= (32'b???????????????????1????????????=>32'b???????????????????0????????????);
		wildcard bins b_1_0_13 	= (32'b??????????????????1?????????????=>32'b??????????????????0?????????????);
		wildcard bins b_1_0_14 	= (32'b?????????????????1??????????????=>32'b?????????????????0??????????????);
		wildcard bins b_1_0_15 	= (32'b????????????????1???????????????=>32'b????????????????0???????????????);
		wildcard bins b_1_0_16 	= (32'b???????????????1????????????????=>32'b???????????????0????????????????);
		wildcard bins b_1_0_17 	= (32'b??????????????1?????????????????=>32'b??????????????0?????????????????);
		wildcard bins b_1_0_18 	= (32'b?????????????1??????????????????=>32'b?????????????0??????????????????);
		wildcard bins b_1_0_19 	= (32'b????????????1???????????????????=>32'b????????????0???????????????????);
		wildcard bins b_1_0_20 	= (32'b???????????1????????????????????=>32'b???????????0????????????????????);
		wildcard bins b_1_0_21 	= (32'b??????????1?????????????????????=>32'b??????????0?????????????????????);
		wildcard bins b_1_0_22 	= (32'b?????????1??????????????????????=>32'b?????????0??????????????????????);
		wildcard bins b_1_0_23 	= (32'b????????1???????????????????????=>32'b????????0???????????????????????);
		wildcard bins b_1_0_24 	= (32'b???????1????????????????????????=>32'b???????0????????????????????????);
		wildcard bins b_1_0_25 	= (32'b??????1?????????????????????????=>32'b??????0?????????????????????????);
		wildcard bins b_1_0_26 	= (32'b?????1??????????????????????????=>32'b?????0??????????????????????????);
		wildcard bins b_1_0_27 	= (32'b????1???????????????????????????=>32'b????0???????????????????????????);
		wildcard bins b_1_0_28 	= (32'b???1????????????????????????????=>32'b???0????????????????????????????);
		wildcard bins b_1_0_29 	= (32'b??1?????????????????????????????=>32'b??0?????????????????????????????);
		wildcard bins b_1_0_30 	= (32'b?1??????????????????????????????=>32'b?0??????????????????????????????);
		wildcard bins b_1_0_31 	= (32'b1???????????????????????????????=>32'b0???????????????????????????????);
		wildcard bins b_0_1_0 	= (32'b???????????????????????????????0=>32'b???????????????????????????????1);
		wildcard bins b_0_1_1 	= (32'b??????????????????????????????0?=>32'b??????????????????????????????1?);
		wildcard bins b_0_1_2 	= (32'b?????????????????????????????0??=>32'b?????????????????????????????1??);
		wildcard bins b_0_1_3 	= (32'b????????????????????????????0???=>32'b????????????????????????????1???);
		wildcard bins b_0_1_4 	= (32'b???????????????????????????0????=>32'b???????????????????????????1????);
		wildcard bins b_0_1_5 	= (32'b??????????????????????????0?????=>32'b??????????????????????????1?????);
		wildcard bins b_0_1_6 	= (32'b?????????????????????????0??????=>32'b?????????????????????????1??????);
		wildcard bins b_0_1_7 	= (32'b????????????????????????0???????=>32'b????????????????????????1???????);
		wildcard bins b_0_1_8 	= (32'b???????????????????????0????????=>32'b???????????????????????1????????);
		wildcard bins b_0_1_9 	= (32'b??????????????????????0?????????=>32'b??????????????????????1?????????);
		wildcard bins b_0_1_10 	= (32'b?????????????????????0??????????=>32'b?????????????????????1??????????);
		wildcard bins b_0_1_11 	= (32'b????????????????????0???????????=>32'b????????????????????1???????????);
		wildcard bins b_0_1_12 	= (32'b???????????????????0????????????=>32'b???????????????????1????????????);
		wildcard bins b_0_1_13 	= (32'b??????????????????0?????????????=>32'b??????????????????1?????????????);
		wildcard bins b_0_1_14 	= (32'b?????????????????0??????????????=>32'b?????????????????1??????????????);
		wildcard bins b_0_1_15 	= (32'b????????????????0???????????????=>32'b????????????????1???????????????);
		wildcard bins b_0_1_16 	= (32'b???????????????0????????????????=>32'b???????????????1????????????????);
		wildcard bins b_0_1_17 	= (32'b??????????????0?????????????????=>32'b??????????????1?????????????????);
		wildcard bins b_0_1_18 	= (32'b?????????????0??????????????????=>32'b?????????????1??????????????????);
		wildcard bins b_0_1_19 	= (32'b????????????0???????????????????=>32'b????????????1???????????????????);
		wildcard bins b_0_1_20 	= (32'b???????????0????????????????????=>32'b???????????1????????????????????);
		wildcard bins b_0_1_21 	= (32'b??????????0?????????????????????=>32'b??????????1?????????????????????);
		wildcard bins b_0_1_22 	= (32'b?????????0??????????????????????=>32'b?????????1??????????????????????);
		wildcard bins b_0_1_23 	= (32'b????????0???????????????????????=>32'b????????1???????????????????????);
		wildcard bins b_0_1_24 	= (32'b???????0????????????????????????=>32'b???????1????????????????????????);
		wildcard bins b_0_1_25 	= (32'b??????0?????????????????????????=>32'b??????1?????????????????????????);
		wildcard bins b_0_1_26 	= (32'b?????0??????????????????????????=>32'b?????1??????????????????????????);
		wildcard bins b_0_1_27 	= (32'b????0???????????????????????????=>32'b????1???????????????????????????);
		wildcard bins b_0_1_28 	= (32'b???0????????????????????????????=>32'b???1????????????????????????????);
		wildcard bins b_0_1_29 	= (32'b??0?????????????????????????????=>32'b??1?????????????????????????????);
		wildcard bins b_0_1_30 	= (32'b?0??????????????????????????????=>32'b?1??????????????????????????????);
		wildcard bins b_0_1_31 	= (32'b0???????????????????????????????=>32'b1???????????????????????????????);
		option.weight = 1;
	 }

	//RS1 special values
	rs1_sp_val: coverpoint unsigned'(rv32i_trans.rs1_val) iff(rv32i_trans.trap==0) {
		bins b0 = {32'b0};
		bins b1 = {32'b00000000000000000000000000000001};
		bins b2 = {32'b11111111111111111111111111111111};
		bins b3 = {32'b01111111111111111111111111111111};
		bins b4 = {32'b10000000000000000000000000000000};
		bins b5 = {32'b10000000000000000000000000000001};
		option.weight = 1;
	 }

	//RS1 value sign
	rs1_val_sign: coverpoint rv32i_trans.rs1_val iff(rv32i_trans.trap==0) {
		bins b0 = {[$:-1]};
		bins b1 = {[1:$]};
		option.weight = 1;
	 }

	//RS2 toggle bits
	rs2_val: coverpoint unsigned'(rv32i_trans.rs2_val) iff(rv32i_trans.trap==0) {
		wildcard bins b_1_0_0 	= (32'b???????????????????????????????1=>32'b???????????????????????????????0);
		wildcard bins b_1_0_1 	= (32'b??????????????????????????????1?=>32'b??????????????????????????????0?);
		wildcard bins b_1_0_2 	= (32'b?????????????????????????????1??=>32'b?????????????????????????????0??);
		wildcard bins b_1_0_3 	= (32'b????????????????????????????1???=>32'b????????????????????????????0???);
		wildcard bins b_1_0_4 	= (32'b???????????????????????????1????=>32'b???????????????????????????0????);
		wildcard bins b_1_0_5 	= (32'b??????????????????????????1?????=>32'b??????????????????????????0?????);
		wildcard bins b_1_0_6 	= (32'b?????????????????????????1??????=>32'b?????????????????????????0??????);
		wildcard bins b_1_0_7 	= (32'b????????????????????????1???????=>32'b????????????????????????0???????);
		wildcard bins b_1_0_8 	= (32'b???????????????????????1????????=>32'b???????????????????????0????????);
		wildcard bins b_1_0_9 	= (32'b??????????????????????1?????????=>32'b??????????????????????0?????????);
		wildcard bins b_1_0_10 	= (32'b?????????????????????1??????????=>32'b?????????????????????0??????????);
		wildcard bins b_1_0_11 	= (32'b????????????????????1???????????=>32'b????????????????????0???????????);
		wildcard bins b_1_0_12 	= (32'b???????????????????1????????????=>32'b???????????????????0????????????);
		wildcard bins b_1_0_13 	= (32'b??????????????????1?????????????=>32'b??????????????????0?????????????);
		wildcard bins b_1_0_14 	= (32'b?????????????????1??????????????=>32'b?????????????????0??????????????);
		wildcard bins b_1_0_15 	= (32'b????????????????1???????????????=>32'b????????????????0???????????????);
		wildcard bins b_1_0_16 	= (32'b???????????????1????????????????=>32'b???????????????0????????????????);
		wildcard bins b_1_0_17 	= (32'b??????????????1?????????????????=>32'b??????????????0?????????????????);
		wildcard bins b_1_0_18 	= (32'b?????????????1??????????????????=>32'b?????????????0??????????????????);
		wildcard bins b_1_0_19 	= (32'b????????????1???????????????????=>32'b????????????0???????????????????);
		wildcard bins b_1_0_20 	= (32'b???????????1????????????????????=>32'b???????????0????????????????????);
		wildcard bins b_1_0_21 	= (32'b??????????1?????????????????????=>32'b??????????0?????????????????????);
		wildcard bins b_1_0_22 	= (32'b?????????1??????????????????????=>32'b?????????0??????????????????????);
		wildcard bins b_1_0_23 	= (32'b????????1???????????????????????=>32'b????????0???????????????????????);
		wildcard bins b_1_0_24 	= (32'b???????1????????????????????????=>32'b???????0????????????????????????);
		wildcard bins b_1_0_25 	= (32'b??????1?????????????????????????=>32'b??????0?????????????????????????);
		wildcard bins b_1_0_26 	= (32'b?????1??????????????????????????=>32'b?????0??????????????????????????);
		wildcard bins b_1_0_27 	= (32'b????1???????????????????????????=>32'b????0???????????????????????????);
		wildcard bins b_1_0_28 	= (32'b???1????????????????????????????=>32'b???0????????????????????????????);
		wildcard bins b_1_0_29 	= (32'b??1?????????????????????????????=>32'b??0?????????????????????????????);
		wildcard bins b_1_0_30 	= (32'b?1??????????????????????????????=>32'b?0??????????????????????????????);
		wildcard bins b_1_0_31 	= (32'b1???????????????????????????????=>32'b0???????????????????????????????);
		wildcard bins b_0_1_0 	= (32'b???????????????????????????????0=>32'b???????????????????????????????1);
		wildcard bins b_0_1_1 	= (32'b??????????????????????????????0?=>32'b??????????????????????????????1?);
		wildcard bins b_0_1_2 	= (32'b?????????????????????????????0??=>32'b?????????????????????????????1??);
		wildcard bins b_0_1_3 	= (32'b????????????????????????????0???=>32'b????????????????????????????1???);
		wildcard bins b_0_1_4 	= (32'b???????????????????????????0????=>32'b???????????????????????????1????);
		wildcard bins b_0_1_5 	= (32'b??????????????????????????0?????=>32'b??????????????????????????1?????);
		wildcard bins b_0_1_6 	= (32'b?????????????????????????0??????=>32'b?????????????????????????1??????);
		wildcard bins b_0_1_7 	= (32'b????????????????????????0???????=>32'b????????????????????????1???????);
		wildcard bins b_0_1_8 	= (32'b???????????????????????0????????=>32'b???????????????????????1????????);
		wildcard bins b_0_1_9 	= (32'b??????????????????????0?????????=>32'b??????????????????????1?????????);
		wildcard bins b_0_1_10 	= (32'b?????????????????????0??????????=>32'b?????????????????????1??????????);
		wildcard bins b_0_1_11 	= (32'b????????????????????0???????????=>32'b????????????????????1???????????);
		wildcard bins b_0_1_12 	= (32'b???????????????????0????????????=>32'b???????????????????1????????????);
		wildcard bins b_0_1_13 	= (32'b??????????????????0?????????????=>32'b??????????????????1?????????????);
		wildcard bins b_0_1_14 	= (32'b?????????????????0??????????????=>32'b?????????????????1??????????????);
		wildcard bins b_0_1_15 	= (32'b????????????????0???????????????=>32'b????????????????1???????????????);
		wildcard bins b_0_1_16 	= (32'b???????????????0????????????????=>32'b???????????????1????????????????);
		wildcard bins b_0_1_17 	= (32'b??????????????0?????????????????=>32'b??????????????1?????????????????);
		wildcard bins b_0_1_18 	= (32'b?????????????0??????????????????=>32'b?????????????1??????????????????);
		wildcard bins b_0_1_19 	= (32'b????????????0???????????????????=>32'b????????????1???????????????????);
		wildcard bins b_0_1_20 	= (32'b???????????0????????????????????=>32'b???????????1????????????????????);
		wildcard bins b_0_1_21 	= (32'b??????????0?????????????????????=>32'b??????????1?????????????????????);
		wildcard bins b_0_1_22 	= (32'b?????????0??????????????????????=>32'b?????????1??????????????????????);
		wildcard bins b_0_1_23 	= (32'b????????0???????????????????????=>32'b????????1???????????????????????);
		wildcard bins b_0_1_24 	= (32'b???????0????????????????????????=>32'b???????1????????????????????????);
		wildcard bins b_0_1_25 	= (32'b??????0?????????????????????????=>32'b??????1?????????????????????????);
		wildcard bins b_0_1_26 	= (32'b?????0??????????????????????????=>32'b?????1??????????????????????????);
		wildcard bins b_0_1_27 	= (32'b????0???????????????????????????=>32'b????1???????????????????????????);
		wildcard bins b_0_1_28 	= (32'b???0????????????????????????????=>32'b???1????????????????????????????);
		wildcard bins b_0_1_29 	= (32'b??0?????????????????????????????=>32'b??1?????????????????????????????);
		wildcard bins b_0_1_30 	= (32'b?0??????????????????????????????=>32'b?1??????????????????????????????);
		wildcard bins b_0_1_31 	= (32'b0???????????????????????????????=>32'b1???????????????????????????????);
		option.weight = 1;
	 }

	//RS2 special values
	rs2_sp_val: coverpoint unsigned'(rv32i_trans.rs2_val) iff(rv32i_trans.trap==0) {
		bins b0 = {32'b0};
		bins b1 = {32'b00000000000000000000000000000001};
		bins b2 = {32'b11111111111111111111111111111111};
		bins b3 = {32'b01111111111111111111111111111111};
		bins b4 = {32'b10000000000000000000000000000000};
		bins b5 = {32'b10000000000000000000000000000001};
		option.weight = 1;
	 }

	//RS2 value sign
	rs2_val_sign: coverpoint rv32i_trans.rs2_val iff(rv32i_trans.trap==0) {
		bins b0 = {[$:-1]};
		bins b1 = {[1:$]};
		option.weight = 1;
	 }

	//12-bit immediate
	imm_12bit: coverpoint unsigned'(rv32i_trans.imm_12bit) iff(rv32i_trans.trap==0) {
		wildcard bins b_1_0_0 	= (12'b???????????1=>12'b???????????0);
		wildcard bins b_1_0_1 	= (12'b??????????1?=>12'b??????????0?);
		wildcard bins b_1_0_2 	= (12'b?????????1??=>12'b?????????0??);
		wildcard bins b_1_0_3 	= (12'b????????1???=>12'b????????0???);
		wildcard bins b_1_0_4 	= (12'b???????1????=>12'b???????0????);
		wildcard bins b_1_0_5 	= (12'b??????1?????=>12'b??????0?????);
		wildcard bins b_1_0_6 	= (12'b?????1??????=>12'b?????0??????);
		wildcard bins b_1_0_7 	= (12'b????1???????=>12'b????0???????);
		wildcard bins b_1_0_8 	= (12'b???1????????=>12'b???0????????);
		wildcard bins b_1_0_9 	= (12'b??1?????????=>12'b??0?????????);
		wildcard bins b_1_0_10 	= (12'b?1??????????=>12'b?0??????????);
		wildcard bins b_1_0_11 	= (12'b1???????????=>12'b0???????????);
		wildcard bins b_0_1_0 	= (12'b???????????0=>12'b???????????1);
		wildcard bins b_0_1_1 	= (12'b??????????0?=>12'b??????????1?);
		wildcard bins b_0_1_2 	= (12'b?????????0??=>12'b?????????1??);
		wildcard bins b_0_1_3 	= (12'b????????0???=>12'b????????1???);
		wildcard bins b_0_1_4 	= (12'b???????0????=>12'b???????1????);
		wildcard bins b_0_1_5 	= (12'b??????0?????=>12'b??????1?????);
		wildcard bins b_0_1_6 	= (12'b?????0??????=>12'b?????1??????);
		wildcard bins b_0_1_7 	= (12'b????0???????=>12'b????1???????);
		wildcard bins b_0_1_8 	= (12'b???0????????=>12'b???1????????);
		wildcard bins b_0_1_9 	= (12'b??0?????????=>12'b??1?????????);
		wildcard bins b_0_1_10 	= (12'b?0??????????=>12'b?1??????????);
		wildcard bins b_0_1_11 	= (12'b0???????????=>12'b1???????????);
		option.weight = 1;
	 }

	//12-bit immediate
	imm_12bit_sign: coverpoint rv32i_trans.imm_12bit iff(rv32i_trans.trap==0) {
		bins b0 = {[$:-1]};
		bins b1 = {0};
		bins b2 = {[1:$]};
		option.weight = 1;
	 }

	//20-bit immediate
	imm_20bit: coverpoint unsigned'(rv32i_trans.imm_20bit) iff(rv32i_trans.trap==0) {
		wildcard bins b_1_0_0 	= (20'b???????????????????1=>20'b???????????????????0);
		wildcard bins b_1_0_1 	= (20'b??????????????????1?=>20'b??????????????????0?);
		wildcard bins b_1_0_2 	= (20'b?????????????????1??=>20'b?????????????????0??);
		wildcard bins b_1_0_3 	= (20'b????????????????1???=>20'b????????????????0???);
		wildcard bins b_1_0_4 	= (20'b???????????????1????=>20'b???????????????0????);
		wildcard bins b_1_0_5 	= (20'b??????????????1?????=>20'b??????????????0?????);
		wildcard bins b_1_0_6 	= (20'b?????????????1??????=>20'b?????????????0??????);
		wildcard bins b_1_0_7 	= (20'b????????????1???????=>20'b????????????0???????);
		wildcard bins b_1_0_8 	= (20'b???????????1????????=>20'b???????????0????????);
		wildcard bins b_1_0_9 	= (20'b??????????1?????????=>20'b??????????0?????????);
		wildcard bins b_1_0_10 	= (20'b?????????1??????????=>20'b?????????0??????????);
		wildcard bins b_1_0_11 	= (20'b????????1???????????=>20'b????????0???????????);
		wildcard bins b_1_0_12 	= (20'b???????1????????????=>20'b???????0????????????);
		wildcard bins b_1_0_13 	= (20'b??????1?????????????=>20'b??????0?????????????);
		wildcard bins b_1_0_14 	= (20'b?????1??????????????=>20'b?????0??????????????);
		wildcard bins b_1_0_15 	= (20'b????1???????????????=>20'b????0???????????????);
		wildcard bins b_1_0_16 	= (20'b???1????????????????=>20'b???0????????????????);
		wildcard bins b_1_0_17 	= (20'b??1?????????????????=>20'b??0?????????????????);
		wildcard bins b_1_0_18 	= (20'b?1??????????????????=>20'b?0??????????????????);
		wildcard bins b_1_0_19 	= (20'b1???????????????????=>20'b0???????????????????);
		wildcard bins b_0_1_0 	= (20'b???????????????????0=>20'b???????????????????1);
		wildcard bins b_0_1_1 	= (20'b??????????????????0?=>20'b??????????????????1?);
		wildcard bins b_0_1_2 	= (20'b?????????????????0??=>20'b?????????????????1??);
		wildcard bins b_0_1_3 	= (20'b????????????????0???=>20'b????????????????1???);
		wildcard bins b_0_1_4 	= (20'b???????????????0????=>20'b???????????????1????);
		wildcard bins b_0_1_5 	= (20'b??????????????0?????=>20'b??????????????1?????);
		wildcard bins b_0_1_6 	= (20'b?????????????0??????=>20'b?????????????1??????);
		wildcard bins b_0_1_7 	= (20'b????????????0???????=>20'b????????????1???????);
		wildcard bins b_0_1_8 	= (20'b???????????0????????=>20'b???????????1????????);
		wildcard bins b_0_1_9 	= (20'b??????????0?????????=>20'b??????????1?????????);
		wildcard bins b_0_1_10 	= (20'b?????????0??????????=>20'b?????????1??????????);
		wildcard bins b_0_1_11 	= (20'b????????0???????????=>20'b????????1???????????);
		wildcard bins b_0_1_12 	= (20'b???????0????????????=>20'b???????1????????????);
		wildcard bins b_0_1_13 	= (20'b??????0?????????????=>20'b??????1?????????????);
		wildcard bins b_0_1_14 	= (20'b?????0??????????????=>20'b?????1??????????????);
		wildcard bins b_0_1_15 	= (20'b????0???????????????=>20'b????1???????????????);
		wildcard bins b_0_1_16 	= (20'b???0????????????????=>20'b???1????????????????);
		wildcard bins b_0_1_17 	= (20'b??0?????????????????=>20'b??1?????????????????);
		wildcard bins b_0_1_18 	= (20'b?0??????????????????=>20'b?1??????????????????);
		wildcard bins b_0_1_19 	= (20'b0???????????????????=>20'b1???????????????????);
		option.weight = 1;
	 }

	//20-bit immediate
	imm_20bit_sign: coverpoint rv32i_trans.imm_20bit iff(rv32i_trans.trap==0) {
		bins b0 = {[$:-1]};
		bins b1 = {0};
		bins b2 = {[1:$]};
		option.weight = 1;
	 }

	// coverpoint for ADD/AND/OR/SUB/XOR
	//war_hazard
	war_hazard_hit: coverpoint rv32i_trans.war_hazard_hit iff(rv32i_trans.trap==0) {
		bins b0 = {1};
		option.weight = 1;
	 }

	//waw_hazard
	waw_hazard_hit: coverpoint rv32i_trans.waw_hazard_hit iff(rv32i_trans.trap==0) {
		bins b0 = {1};
		option.weight = 1;
	 }

	//raw_hazard
	raw_hazard_hit: coverpoint rv32i_trans.raw_hazard_hit iff(rv32i_trans.trap==0) {
		bins b0 = {1};
		option.weight = 1;
	 }

	// coverpoint for SLLI/SRLI/SRAL
	//immediate values used by shift instruction
	imm_shift: coverpoint rv32i_trans.imm_12bit iff(rv32i_trans.trap==0) {
		bins b0 = {[0:5]};
		bins b1 = {[6:10]};
		bins b2 = {[11:15]};
		bins b3 = {[16:20]};
		bins b4 = {[21:25]};
		bins b5 = {[26:30]};
		bins b6 = {31};
		option.weight = 1;
	 }

	// coverpoint for BEQ/BNE/BLT/BGE/BLTU/BGEU
	//rs1_val == rs2_val
	rs1_val_eq_rs2_val: coverpoint rv32i_trans.rs1_val==rv32i_trans.rs2_val iff(rv32i_trans.trap==0) {
		bins b0 = {0};
		bins b1 = {1};
		option.weight = 1;
	 }

	// coverpoint for LH/LHU/LW/SH/SW
	//Unaligned memory address when load/store 2 bytes
	half_word_mem_unalign: coverpoint (rv32i_trans.rs1_val+rv32i_trans.imm_12bit)%2 iff(rv32i_trans.trap==0) {
		bins b0 = {0};
		bins b1 = {1};
		option.weight = 1;
	 }

	//Unaligned memory address when load/store 4 bytes
	word_mem_unalign: coverpoint (rv32i_trans.rs1_val+rv32i_trans.imm_12bit)%4 iff(rv32i_trans.trap==0) {
		bins b0 = {0};
		bins b1 = {1};
		bins b2 = {2};
		bins b3 = {3};
		option.weight = 1;
	 }

	//Unaligned memory address when load/store 4 bytes
	mem_start_addr: coverpoint (rv32i_trans.rs1_val+rv32i_trans.imm_12bit)%16 iff(rv32i_trans.trap==0) {
		bins b0 = {0};
		bins b1 = {1};
		bins b2 = {2};
		bins b3 = {3};
		bins b4 = {4};
		bins b5 = {5};
		bins b6 = {6};
		bins b7 = {7};
		bins b8 = {8};
		bins b9 = {9};
		bins b10 = {10};
		bins b11 = {11};
		bins b12 = {12};
		bins b13 = {13};
		bins b14 = {14};
		bins b15 = {15};
		option.weight = 1;
	 }

	// coverpoint for jal/lui/auipc
	//20-bit immediate is 0
	imm_zero: coverpoint unsigned'(rv32i_trans.imm_20bit) iff(rv32i_trans.trap==0) {
		bins b0 = {0};
		option.weight = 1;
	 }

	// coverpoint for fence
	//4'b0000:normal fence
	//4'b1000:fence rw.rw
	fm: coverpoint rv32i_trans.fm iff(rv32i_trans.trap==0) {
		bins b0 = {4'b0000};
		bins b1 = {4'b1000};
		option.weight = 1;
	 }

	//predecessors,
	//Bit3:Input,bit2:output,bit3:read,bit0:write
	pred: coverpoint rv32i_trans.pred iff(rv32i_trans.trap==0) {
		bins b0 = {4'b0000};
		bins b1 = {4'b0001};
		bins b2 = {4'b0010};
		bins b3 = {4'b0011};
		bins b4 = {4'b0100};
		bins b5 = {4'b0101};
		bins b6 = {4'b0110};
		bins b7 = {4'b0111};
		bins b8 = {4'b1000};
		bins b9 = {4'b1001};
		bins b10 = {4'b1010};
		bins b11 = {4'b1011};
		bins b12 = {4'b1100};
		bins b13 = {4'b1101};
		bins b14 = {4'b1110};
		bins b15 = {4'b1111};
		option.weight = 1;
	 }

	//Successors,
	//Bit3:Input,bit2:output,bit3:read,bit0:write
	succ: coverpoint rv32i_trans.succ iff(rv32i_trans.trap==0) {
		bins b0 = {4'b0000};
		bins b1 = {4'b0001};
		bins b2 = {4'b0010};
		bins b3 = {4'b0011};
		bins b4 = {4'b0100};
		bins b5 = {4'b0101};
		bins b6 = {4'b0110};
		bins b7 = {4'b0111};
		bins b8 = {4'b1000};
		bins b9 = {4'b1001};
		bins b10 = {4'b1010};
		bins b11 = {4'b1011};
		bins b12 = {4'b1100};
		bins b13 = {4'b1101};
		bins b14 = {4'b1110};
		bins b15 = {4'b1111};
		option.weight = 1;
	 }

	// base cross
	//Cross ADD instruction  and register assignment
	cr_add_rs1_rs2_rd: cross add,rs1_addr,rs2_addr,rd_addr {
		option.weight = 1;
	}

	//Cross ADD instruction  and RS1 toggle bits
	cr_add_rs1_val: cross add,rs1_val {
		option.weight = 1;
	}

	//Cross ADD instruction  and RS1 special values
	cr_add_rs1_sp_val: cross add,rs1_sp_val {
		option.weight = 1;
	}

	//Cross ADD instruction  and RS1 value sign
	cr_add_rs1_val_sign: cross add,rs1_val_sign {
		option.weight = 1;
	}

	//Cross ADD instruction  and RS2 toggle bits
	cr_add_rs2_val: cross add,rs2_val {
		option.weight = 1;
	}

	//Cross ADD instruction  and RS2 special values
	cr_add_rs2_sp_val: cross add,rs2_sp_val {
		option.weight = 1;
	}

	//Cross ADD instruction  and RS2 value sign
	cr_add_rs2_val_sign: cross add,rs2_val_sign {
		option.weight = 1;
	}

	//Cross ADD instruction  and RD toggle bits
	cr_add_rd_val: cross add,rd_val {
		option.weight = 1;
	}

	//Cross ADD instruction  and RD special values
	cr_add_rd_sp_val: cross add,rd_sp_val {
		option.weight = 1;
	}

	//Cross ADD instruction  and RD value sign
	cr_add_rd_val_sign: cross add,rd_val_sign {
		option.weight = 1;
	}

	//Cross ADD instruction  and WAR hazard
	cr_add_war_hazard: cross add,war_hazard_hit {
		option.weight = 1;
	}

	//Cross ADD instruction  and WAW hazard
	cr_add_waw_hazard: cross add,waw_hazard_hit {
		option.weight = 1;
	}

	//Cross ADD instruction  and RAW hazard
	cr_add_raw_hazard: cross add,raw_hazard_hit {
		option.weight = 1;
	}

	//Cross SUB instruction  and register assignment
	cr_sub_rs1_rs2_rd: cross sub,rs1_addr,rs2_addr,rd_addr {
		option.weight = 1;
	}

	//Cross SUB instruction  and RS1 toggle bits
	cr_sub_rs1_val: cross sub,rs1_val {
		option.weight = 1;
	}

	//Cross SUB instruction  and RS1 special values
	cr_sub_rs1_sp_val: cross sub,rs1_sp_val {
		option.weight = 1;
	}

	//Cross SUB instruction  and RS1 value sign
	cr_sub_rs1_val_sign: cross sub,rs1_val_sign {
		option.weight = 1;
	}

	//Cross SUB instruction  and RS2 toggle bits
	cr_sub_rs2_val: cross sub,rs2_val {
		option.weight = 1;
	}

	//Cross SUB instruction  and RS2 special values
	cr_sub_rs2_sp_val: cross sub,rs2_sp_val {
		option.weight = 1;
	}

	//Cross SUB instruction  and RS2 value sign
	cr_sub_rs2_val_sign: cross sub,rs2_val_sign {
		option.weight = 1;
	}

	//Cross SUB instruction  and RD toggle bits
	cr_sub_rd_val: cross sub,rd_val {
		option.weight = 1;
	}

	//Cross SUB instruction  and RD special values
	cr_sub_rd_sp_val: cross sub,rd_sp_val {
		option.weight = 1;
	}

	//Cross SUB instruction  and RD value sign
	cr_sub_rd_val_sign: cross sub,rd_val_sign {
		option.weight = 1;
	}

	//Cross SUB instruction  and WAR hazard
	cr_sub_war_hazard: cross sub,war_hazard_hit {
		option.weight = 1;
	}

	//Cross SUB instruction  and WAW hazard
	cr_sub_waw_hazard: cross sub,waw_hazard_hit {
		option.weight = 1;
	}

	//Cross SUB instruction  and RAW hazard
	cr_sub_raw_hazard: cross sub,raw_hazard_hit {
		option.weight = 1;
	}

	//Cross XOR instruction  and register assignment
	cr_xor_rs1_rs2_rd: cross cp_xor,rs1_addr,rs2_addr,rd_addr {
		option.weight = 1;
	}

	//Cross XOR instruction  and RS1 toggle bits
	cr_xor_rs1_val: cross cp_xor,rs1_val {
		option.weight = 1;
	}

	//Cross XOR instruction  and RS1 special values
	cr_xor_rs1_sp_val: cross cp_xor,rs1_sp_val {
		option.weight = 1;
	}

	//Cross XOR instruction  and RS1 value sign
	cr_xor_rs1_val_sign: cross cp_xor,rs1_val_sign {
		option.weight = 1;
	}

	//Cross XOR instruction  and RS2 toggle bits
	cr_xor_rs2_val: cross cp_xor,rs2_val {
		option.weight = 1;
	}

	//Cross XOR instruction  and RS2 special values
	cr_xor_rs2_sp_val: cross cp_xor,rs2_sp_val {
		option.weight = 1;
	}

	//Cross XOR instruction  and RS2 value sign
	cr_xor_rs2_val_sign: cross cp_xor,rs2_val_sign {
		option.weight = 1;
	}

	//Cross XOR instruction  and RD toggle bits
	cr_xor_rd_val: cross cp_xor,rd_val {
		option.weight = 1;
	}

	//Cross XOR instruction  and RD special values
	cr_xor_rd_sp_val: cross cp_xor,rd_sp_val {
		option.weight = 1;
	}

	//Cross XOR instruction  and RD value sign
	cr_xor_rd_val_sign: cross cp_xor,rd_val_sign {
		option.weight = 1;
	}

	//Cross XOR instruction  and WAR hazard
	cr_xor_war_hazard: cross cp_xor,war_hazard_hit {
		option.weight = 1;
	}

	//Cross XOR instruction  and WAW hazard
	cr_xor_waw_hazard: cross cp_xor,waw_hazard_hit {
		option.weight = 1;
	}

	//Cross XOR instruction  and RAW hazard
	cr_xor_raw_hazard: cross cp_xor,raw_hazard_hit {
		option.weight = 1;
	}

	//Cross OR instruction  and register assignment
	cr_or_rs1_rs2_rd: cross cp_or,rs1_addr,rs2_addr,rd_addr {
		option.weight = 1;
	}

	//Cross OR instruction  and RS1 toggle bits
	cr_or_rs1_val: cross cp_or,rs1_val {
		option.weight = 1;
	}

	//Cross OR instruction  and RS1 special values
	cr_or_rs1_sp_val: cross cp_or,rs1_sp_val {
		option.weight = 1;
	}

	//Cross OR instruction  and RS1 value sign
	cr_or_rs1_val_sign: cross cp_or,rs1_val_sign {
		option.weight = 1;
	}

	//Cross OR instruction  and RS2 toggle bits
	cr_or_rs2_val: cross cp_or,rs2_val {
		option.weight = 1;
	}

	//Cross OR instruction  and RS2 special values
	cr_or_rs2_sp_val: cross cp_or,rs2_sp_val {
		option.weight = 1;
	}

	//Cross OR instruction  and RS2 value sign
	cr_or_rs2_val_sign: cross cp_or,rs2_val_sign {
		option.weight = 1;
	}

	//Cross OR instruction  and RD toggle bits
	cr_or_rd_val: cross cp_or,rd_val {
		option.weight = 1;
	}

	//Cross OR instruction  and RD special values
	cr_or_rd_sp_val: cross cp_or,rd_sp_val {
		option.weight = 1;
	}

	//Cross OR instruction  and RD value sign
	cr_or_rd_val_sign: cross cp_or,rd_val_sign {
		option.weight = 1;
	}

	//Cross OR instruction  and WAR hazard
	cr_or_war_hazard: cross cp_or,war_hazard_hit {
		option.weight = 1;
	}

	//Cross OR instruction  and WAW hazard
	cr_or_waw_hazard: cross cp_or,waw_hazard_hit {
		option.weight = 1;
	}

	//Cross OR instruction  and RAW hazard
	cr_or_raw_hazard: cross cp_or,raw_hazard_hit {
		option.weight = 1;
	}

	//Cross AND instruction  and register assignment
	cr_and_rs1_rs2_rd: cross cp_and,rs1_addr,rs2_addr,rd_addr {
		option.weight = 1;
	}

	//Cross AND instruction  and RS1 toggle bits
	cr_and_rs1_val: cross cp_and,rs1_val {
		option.weight = 1;
	}

	//Cross AND instruction  and RS1 special values
	cr_and_rs1_sp_val: cross cp_and,rs1_sp_val {
		option.weight = 1;
	}

	//Cross AND instruction  and RS1 value sign
	cr_and_rs1_val_sign: cross cp_and,rs1_val_sign {
		option.weight = 1;
	}

	//Cross AND instruction  and RS2 toggle bits
	cr_and_rs2_val: cross cp_and,rs2_val {
		option.weight = 1;
	}

	//Cross AND instruction  and RS2 special values
	cr_and_rs2_sp_val: cross cp_and,rs2_sp_val {
		option.weight = 1;
	}

	//Cross AND instruction  and RS2 value sign
	cr_and_rs2_val_sign: cross cp_and,rs2_val_sign {
		option.weight = 1;
	}

	//Cross AND instruction  and RD toggle bits
	cr_and_rd_val: cross cp_and,rd_val {
		option.weight = 1;
	}

	//Cross AND instruction  and RD special values
	cr_and_rd_sp_val: cross cp_and,rd_sp_val {
		option.weight = 1;
	}

	//Cross AND instruction  and RD value sign
	cr_and_rd_val_sign: cross cp_and,rd_val_sign {
		option.weight = 1;
	}

	//Cross AND instruction  and WAR hazard
	cr_and_war_hazard: cross cp_and,war_hazard_hit {
		option.weight = 1;
	}

	//Cross AND instruction  and WAW hazard
	cr_and_waw_hazard: cross cp_and,waw_hazard_hit {
		option.weight = 1;
	}

	//Cross AND instruction  and RAW hazard
	cr_and_raw_hazard: cross cp_and,raw_hazard_hit {
		option.weight = 1;
	}

	//Cross SLL instruction  and register assignment
	cr_sll_rs1_rs2_rd: cross sll,rs1_addr,rs2_addr,rd_addr {
		option.weight = 1;
	}

	//Cross SLL instruction  and RS1 toggle bits
	cr_sll_rs1_val: cross sll,rs1_val {
		option.weight = 1;
	}

	//Cross SLL instruction  and RS1 special values
	cr_sll_rs1_sp_val: cross sll,rs1_sp_val {
		option.weight = 1;
	}

	//Cross SLL instruction  and RS1 value sign
	cr_sll_rs1_val_sign: cross sll,rs1_val_sign {
		option.weight = 1;
	}

	//Cross SLL instruction  and RS2 toggle bits
	cr_sll_rs2_val: cross sll,rs2_val {
		option.weight = 1;
	}

	//Cross SLL instruction  and RS2 special values
	cr_sll_rs2_sp_val: cross sll,rs2_sp_val {
		option.weight = 1;
	}

	//Cross SLL instruction  and RS2 value sign
	cr_sll_rs2_val_sign: cross sll,rs2_val_sign {
		option.weight = 1;
	}

	//Cross SLL instruction  and RD toggle bits
	cr_sll_rd_val: cross sll,rd_val {
		option.weight = 1;
	}

	//Cross SLL instruction  and RD special values
	cr_sll_rd_sp_val: cross sll,rd_sp_val {
		option.weight = 1;
	}

	//Cross SLL instruction  and RD value sign
	cr_sll_rd_val_sign: cross sll,rd_val_sign {
		option.weight = 1;
	}

	//Cross SRL instruction  and register assignment
	cr_srl_rs1_rs2_rd: cross srl,rs1_addr,rs2_addr,rd_addr {
		option.weight = 1;
	}

	//Cross SRL instruction  and RS1 toggle bits
	cr_srl_rs1_val: cross srl,rs1_val {
		option.weight = 1;
	}

	//Cross SRL instruction  and RS1 special values
	cr_srl_rs1_sp_val: cross srl,rs1_sp_val {
		option.weight = 1;
	}

	//Cross SRL instruction  and RS1 value sign
	cr_srl_rs1_val_sign: cross srl,rs1_val_sign {
		option.weight = 1;
	}

	//Cross SRL instruction  and RS2 toggle bits
	cr_srl_rs2_val: cross srl,rs2_val {
		option.weight = 1;
	}

	//Cross SRL instruction  and RS2 special values
	cr_srl_rs2_sp_val: cross srl,rs2_sp_val {
		option.weight = 1;
	}

	//Cross SRL instruction  and RS2 value sign
	cr_srl_rs2_val_sign: cross srl,rs2_val_sign {
		option.weight = 1;
	}

	//Cross SRL instruction  and RD toggle bits
	cr_srl_rd_val: cross srl,rd_val {
		option.weight = 1;
	}

	//Cross SRL instruction  and RD special values
	cr_srl_rd_sp_val: cross srl,rd_sp_val {
		option.weight = 1;
	}

	//Cross SRL instruction  and RD value sign
	cr_srl_rd_val_sign: cross srl,rd_val_sign {
		option.weight = 1;
	}

	//Cross SRA instruction  and register assignment
	cr_sra_rs1_rs2_rd: cross sra,rs1_addr,rs2_addr,rd_addr {
		option.weight = 1;
	}

	//Cross SRA instruction  and RS1 toggle bits
	cr_sra_rs1_val: cross sra,rs1_val {
		option.weight = 1;
	}

	//Cross SRA instruction  and RS1 special values
	cr_sra_rs1_sp_val: cross sra,rs1_sp_val {
		option.weight = 1;
	}

	//Cross SRA instruction  and RS1 value sign
	cr_sra_rs1_val_sign: cross sra,rs1_val_sign {
		option.weight = 1;
	}

	//Cross SRA instruction  and RS2 toggle bits
	cr_sra_rs2_val: cross sra,rs2_val {
		option.weight = 1;
	}

	//Cross SRA instruction  and RS2 special values
	cr_sra_rs2_sp_val: cross sra,rs2_sp_val {
		option.weight = 1;
	}

	//Cross SRA instruction  and RS2 value sign
	cr_sra_rs2_val_sign: cross sra,rs2_val_sign {
		option.weight = 1;
	}

	//Cross SRA instruction  and RD toggle bits
	cr_sra_rd_val: cross sra,rd_val {
		option.weight = 1;
	}

	//Cross SRA instruction  and RD special values
	cr_sra_rd_sp_val: cross sra,rd_sp_val {
		option.weight = 1;
	}

	//Cross SRA instruction  and RD value sign
	cr_sra_rd_val_sign: cross sra,rd_val_sign {
		option.weight = 1;
	}

	//Cross SLT instruction  and register assignment
	cr_slt_rs1_rs2_rd: cross slt,rs1_addr,rs2_addr,rd_addr {
		option.weight = 1;
	}

	//Cross SLT instruction  and RS1 toggle bits
	cr_slt_rs1_val: cross slt,rs1_val {
		option.weight = 1;
	}

	//Cross SLT instruction  and RS1 special values
	cr_slt_rs1_sp_val: cross slt,rs1_sp_val {
		option.weight = 1;
	}

	//Cross SLT instruction  and RS1 value sign
	cr_slt_rs1_val_sign: cross slt,rs1_val_sign {
		option.weight = 1;
	}

	//Cross SLT instruction  and RS2 toggle bits
	cr_slt_rs2_val: cross slt,rs2_val {
		option.weight = 1;
	}

	//Cross SLT instruction  and RS2 special values
	cr_slt_rs2_sp_val: cross slt,rs2_sp_val {
		option.weight = 1;
	}

	//Cross SLT instruction  and RS2 value sign
	cr_slt_rs2_val_sign: cross slt,rs2_val_sign {
		option.weight = 1;
	}

	//Cross SLT instruction  and RD toggle bits
	cr_slt_rd_val: cross slt,rd_val {
		option.weight = 1;
	}

	//Cross SLT instruction  and RD special values
	cr_slt_rd_sp_val: cross slt,rd_sp_val {
		option.weight = 1;
	}

	//Cross SLT instruction  and RD value sign
	cr_slt_rd_val_sign: cross slt,rd_val_sign {
		option.weight = 1;
	}

	//Cross SLTU instruction  and register assignment
	cr_sltu_rs1_rs2_rd: cross sltu,rs1_addr,rs2_addr,rd_addr {
		option.weight = 1;
	}

	//Cross SLTU instruction  and RS1 toggle bits
	cr_sltu_rs1_val: cross sltu,rs1_val {
		option.weight = 1;
	}

	//Cross SLTU instruction  and RS1 special values
	cr_sltu_rs1_sp_val: cross sltu,rs1_sp_val {
		option.weight = 1;
	}

	//Cross SLTU instruction  and RS2 toggle bits
	cr_sltu_rs2_val: cross sltu,rs2_val {
		option.weight = 1;
	}

	//Cross SLTU instruction  and RS2 special values
	cr_sltu_rs2_sp_val: cross sltu,rs2_sp_val {
		option.weight = 1;
	}

	//Cross SLTU instruction  and RD toggle bits
	cr_sltu_rd_val: cross sltu,rd_val {
		option.weight = 1;
	}

	//Cross SLTU instruction  and RD special values
	cr_sltu_rd_sp_val: cross sltu,rd_sp_val {
		option.weight = 1;
	}

	//Cross ADDI instruction  and register assignment
	cr_addi_rs1_rd: cross addi,rs1_addr,rd_addr {
		option.weight = 1;
	}

	//Cross ADDI instruction  and RS1 toggle bits
	cr_addi_rs1_val: cross addi,rs1_val {
		option.weight = 1;
	}

	//Cross ADDI instruction  and RS1 special values
	cr_addi_rs1_sp_val: cross addi,rs1_sp_val {
		option.weight = 1;
	}

	//Cross ADDI instruction  and RS1 value sign
	cr_addi_rs1_val_sign: cross addi,rs1_val_sign {
		option.weight = 1;
	}

	//Cross ADDI instruction  and immediate toggle bits
	cr_addi_imm: cross addi,imm_12bit {
		option.weight = 1;
	}

	//Cross ADDI instruction  and immediate value sign
	cr_addi_imm_sign: cross addi,imm_12bit_sign {
		option.weight = 1;
	}

	//Cross ADDI instruction  and RD toggle bits
	cr_addi_rd_val: cross addi,rd_val {
		option.weight = 1;
	}

	//Cross ADDI instruction  and RD special values
	cr_addi_rd_sp_val: cross addi,rd_sp_val {
		option.weight = 1;
	}

	//Cross ADDI instruction  and RD value sign
	cr_addi_rd_val_sign: cross addi,rd_val_sign {
		option.weight = 1;
	}

	//Cross XORI instruction  and register assignment
	cr_xori_rs1_rd: cross xori,rs1_addr,rd_addr {
		option.weight = 1;
	}

	//Cross XORI instruction  and RS1 toggle bits
	cr_xori_rs1_val: cross xori,rs1_val {
		option.weight = 1;
	}

	//Cross XORI instruction  and RS1 special values
	cr_xori_rs1_sp_val: cross xori,rs1_sp_val {
		option.weight = 1;
	}

	//Cross XORI instruction  and RS1 value sign
	cr_xori_rs1_val_sign: cross xori,rs1_val_sign {
		option.weight = 1;
	}

	//Cross XORI instruction  and immediate toggle bits
	cr_xori_imm: cross xori,imm_12bit {
		option.weight = 1;
	}

	//Cross XORI instruction  and immediate value sign
	cr_xori_imm_sign: cross xori,imm_12bit_sign {
		option.weight = 1;
	}

	//Cross XORI instruction  and RD toggle bits
	cr_xori_rd_val: cross xori,rd_val {
		option.weight = 1;
	}

	//Cross XORI instruction  and RD special values
	cr_xori_rd_sp_val: cross xori,rd_sp_val {
		option.weight = 1;
	}

	//Cross XORI instruction  and RD value sign
	cr_xori_rd_val_sign: cross xori,rd_val_sign {
		option.weight = 1;
	}

	//Cross ORI instruction  and register assignment
	cr_ori_rs1_rd: cross ori,rs1_addr,rd_addr {
		option.weight = 1;
	}

	//Cross ORI instruction  and RS1 toggle bits
	cr_ori_rs1_val: cross ori,rs1_val {
		option.weight = 1;
	}

	//Cross ORI instruction  and RS1 special values
	cr_ori_rs1_sp_val: cross ori,rs1_sp_val {
		option.weight = 1;
	}

	//Cross ORI instruction  and RS1 value sign
	cr_ori_rs1_val_sign: cross ori,rs1_val_sign {
		option.weight = 1;
	}

	//Cross ORI instruction  and immediate toggle bits
	cr_ori_imm: cross ori,imm_12bit {
		option.weight = 1;
	}

	//Cross ORI instruction  and immediate value sign
	cr_ori_imm_sign: cross ori,imm_12bit_sign {
		option.weight = 1;
	}

	//Cross ORI instruction  and RD toggle bits
	cr_ori_rd_val: cross ori,rd_val {
		option.weight = 1;
	}

	//Cross ORI instruction  and RD special values
	cr_ori_rd_sp_val: cross ori,rd_sp_val {
		option.weight = 1;
	}

	//Cross ORI instruction  and RD value sign
	cr_ori_rd_val_sign: cross ori,rd_val_sign {
		option.weight = 1;
	}

	//Cross ANDI instruction  and register assignment
	cr_andi_rs1_rd: cross andi,rs1_addr,rd_addr {
		option.weight = 1;
	}

	//Cross ANDI instruction  and RS1 toggle bits
	cr_andi_rs1_val: cross andi,rs1_val {
		option.weight = 1;
	}

	//Cross ANDI instruction  and RS1 special values
	cr_andi_rs1_sp_val: cross andi,rs1_sp_val {
		option.weight = 1;
	}

	//Cross ANDI instruction  and RS1 value sign
	cr_andi_rs1_val_sign: cross andi,rs1_val_sign {
		option.weight = 1;
	}

	//Cross ANDI instruction  and immediate toggle bits
	cr_andi_imm: cross andi,imm_12bit {
		option.weight = 1;
	}

	//Cross ANDI instruction  and immediate value sign
	cr_andi_imm_sign: cross andi,imm_12bit_sign {
		option.weight = 1;
	}

	//Cross ANDI instruction  and RD toggle bits
	cr_andi_rd_val: cross andi,rd_val {
		option.weight = 1;
	}

	//Cross ANDI instruction  and RD special values
	cr_andi_rd_sp_val: cross andi,rd_sp_val {
		option.weight = 1;
	}

	//Cross ANDI instruction  and RD value sign
	cr_andi_rd_val_sign: cross andi,rd_val_sign {
		option.weight = 1;
	}

	//Cross SLLI instruction  and register assignment
	cr_slli_rs1_rd: cross slli,rs1_addr,rd_addr {
		option.weight = 1;
	}

	//Cross SLLI instruction  and RS1 toggle bits
	cr_slli_rs1_val: cross slli,rs1_val {
		option.weight = 1;
	}

	//Cross SLLI instruction  and RS1 special values
	cr_slli_rs1_sp_val: cross slli,rs1_sp_val {
		option.weight = 1;
	}

	//Cross SLLI instruction  and RS1 value sign
	cr_slli_rs1_val_sign: cross slli,rs1_val_sign {
		option.weight = 1;
	}

	//Cross SLLI instruction  and immediate toggle bits
	cr_slli_imm: cross slli,imm_shift {
		option.weight = 1;
	}

	//Cross SLLI instruction  and RD toggle bits
	cr_slli_rd_val: cross slli,rd_val {
		option.weight = 1;
	}

	//Cross SLLI instruction  and RD special values
	cr_slli_rd_sp_val: cross slli,rd_sp_val {
		option.weight = 1;
	}

	//Cross SLLI instruction  and RD value sign
	cr_slli_rd_val_sign: cross slli,rd_val_sign {
		option.weight = 1;
	}

	//Cross SRLI instruction  and register assignment
	cr_srli_rs1_rd: cross srli,rs1_addr,rd_addr {
		option.weight = 1;
	}

	//Cross SRLI instruction  and RS1 toggle bits
	cr_srli_rs1_val: cross srli,rs1_val {
		option.weight = 1;
	}

	//Cross SRLI instruction  and RS1 special values
	cr_srli_rs1_sp_val: cross srli,rs1_sp_val {
		option.weight = 1;
	}

	//Cross SRLI instruction  and RS1 value sign
	cr_srli_rs1_val_sign: cross srli,rs1_val_sign {
		option.weight = 1;
	}

	//Cross SRLI instruction  and immediate toggle bits
	cr_srli_imm: cross srli,imm_shift {
		option.weight = 1;
	}

	//Cross SRLI instruction  and RD toggle bits
	cr_srli_rd_val: cross srli,rd_val {
		option.weight = 1;
	}

	//Cross SRLI instruction  and RD special values
	cr_srli_rd_sp_val: cross srli,rd_sp_val {
		option.weight = 1;
	}

	//Cross SRLI instruction  and RD value sign
	cr_srli_rd_val_sign: cross srli,rd_val_sign {
		option.weight = 1;
	}

	//Cross SRAI instruction  and register assignment
	cr_srai_rs1_rd: cross srai,rs1_addr,rd_addr {
		option.weight = 1;
	}

	//Cross SRAI instruction  and RS1 toggle bits
	cr_srai_rs1_val: cross srai,rs1_val {
		option.weight = 1;
	}

	//Cross SRAI instruction  and RS1 special values
	cr_srai_rs1_sp_val: cross srai,rs1_sp_val {
		option.weight = 1;
	}

	//Cross SRAI instruction  and RS1 value sign
	cr_srai_rs1_val_sign: cross srai,rs1_val_sign {
		option.weight = 1;
	}

	//Cross SRAI instruction  and immediate toggle bits
	cr_srai_imm: cross srai,imm_shift {
		option.weight = 1;
	}

	//Cross SRAI instruction  and RD toggle bits
	cr_srai_rd_val: cross srai,rd_val {
		option.weight = 1;
	}

	//Cross SRAI instruction  and RD special values
	cr_srai_rd_sp_val: cross srai,rd_sp_val {
		option.weight = 1;
	}

	//Cross SRAI instruction  and RD value sign
	cr_srai_rd_val_sign: cross srai,rd_val_sign {
		option.weight = 1;
	}

	//Cross SLTI instruction  and register assignment
	cr_slti_rs1_rd: cross slti,rs1_addr,rd_addr {
		option.weight = 1;
	}

	//Cross SLTI instruction  and RS1 toggle bits
	cr_slti_rs1_val: cross slti,rs1_val {
		option.weight = 1;
	}

	//Cross SLTI instruction  and RS1 special values
	cr_slti_rs1_sp_val: cross slti,rs1_sp_val {
		option.weight = 1;
	}

	//Cross SLTI instruction  and RS1 value sign
	cr_slti_rs1_val_sign: cross slti,rs1_val_sign {
		option.weight = 1;
	}

	//Cross SLTI instruction  and immediate toggle bits
	cr_slti_imm: cross slti,imm_12bit {
		option.weight = 1;
	}

	//Cross SLTI instruction  and immediate value sign
	cr_slti_imm_sign: cross slti,imm_12bit_sign {
		option.weight = 1;
	}

	//Cross SLTI instruction  and RD toggle bits
	cr_slti_rd_val: cross slti,rd_val {
		option.weight = 1;
	}

	//Cross SLTI instruction  and RD special values
	cr_slti_rd_sp_val: cross slti,rd_sp_val {
		option.weight = 1;
	}

	//Cross SLTI instruction  and RD value sign
	cr_slti_rd_val_sign: cross slti,rd_val_sign {
		option.weight = 1;
	}

	//Cross SLTIU instruction  and register assignment
	cr_sltiu_rs1_rd: cross sltiu,rs1_addr,rd_addr {
		option.weight = 1;
	}

	//Cross SLTIU instruction  and RS1 toggle bits
	cr_sltiu_rs1_val: cross sltiu,rs1_val {
		option.weight = 1;
	}

	//Cross SLTIU instruction  and RS1 special values
	cr_sltiu_rs1_sp_val: cross sltiu,rs1_sp_val {
		option.weight = 1;
	}

	//Cross SLTIU instruction  and immediate toggle bits
	cr_sltiu_imm: cross sltiu,imm_12bit {
		option.weight = 1;
	}

	//Cross SLTIU instruction  and RD toggle bits
	cr_sltiu_rd_val: cross sltiu,rd_val {
		option.weight = 1;
	}

	//Cross SLTIU instruction  and RD special values
	cr_sltiu_rd_sp_val: cross sltiu,rd_sp_val {
		option.weight = 1;
	}

	//Cross LB instruction  and RD  assignment
	cr_lb_rd: cross lb,rd_addr {
		option.weight = 1;
	}

	//Cross LB instruction  and RS1 assignment
	cr_lb_rs1: cross lb,rs1_addr {
		option.weight = 1;
	}

	//Cross LB instruction  and immediate toggle bits
	cr_lb_imm: cross lb,imm_12bit {
		option.weight = 1;
	}

	//Cross LB instruction  and immediate value sign
	cr_lb_imm_sign: cross lb,imm_12bit_sign {
		option.weight = 1;
	}

	//Cross LB instruction  and RD toggle bits
	cr_lb_rd_val: cross lb,rd_val {
		option.weight = 1;
	}

	//Cross LB instruction  and RD special values
	cr_lb_rd_sp_val: cross lb,rd_sp_val {
		option.weight = 1;
	}

	//Cross LH instruction  and RD  assignment
	cr_lh_rd: cross lh,rd_addr {
		option.weight = 1;
	}

	//Cross LH instruction  and RS1 assignment
	cr_lh_rs1: cross lh,rs1_addr {
		option.weight = 1;
	}

	//Cross LH instruction  and immediate toggle bits
	cr_lh_imm: cross lh,imm_12bit {
		option.weight = 1;
	}

	//Cross LH instruction  and immediate value sign
	cr_lh_imm_sign: cross lh,imm_12bit_sign {
		option.weight = 1;
	}

	//Cross LH instruction  and RD toggle bits
	cr_lh_rd_val: cross lh,rd_val {
		option.weight = 1;
	}

	//Cross LH instruction  and RD special values
	cr_lh_rd_sp_val: cross lh,rd_sp_val {
		option.weight = 1;
	}

	//Cross LH instruction  and aligned/misaligned memory address
	cr_lh_mem_unalign: cross lh,half_word_mem_unalign {
		option.weight = 1;
	}

	//Cross LH instruction  and aligned/misaligned memory address
	cr_lh_mem_start_addr: cross lh,mem_start_addr {
		option.weight = 1;
	}

	//Cross LW instruction  and RD  assignment
	cr_lw_rd: cross lw,rd_addr {
		option.weight = 1;
	}

	//Cross LW instruction  and RS1 assignment
	cr_lw_rs1: cross lw,rs1_addr {
		option.weight = 1;
	}

	//Cross LW instruction  and immediate toggle bits
	cr_lw_imm: cross lw,imm_12bit {
		option.weight = 1;
	}

	//Cross LW instruction  and immediate value sign
	cr_lw_imm_sign: cross lw,imm_12bit_sign {
		option.weight = 1;
	}

	//Cross LW instruction  and RD toggle bits
	cr_lw_rd_val: cross lw,rd_val {
		option.weight = 1;
	}

	//Cross LW instruction  and RD special values
	cr_lw_rd_sp_val: cross lw,rd_sp_val {
		option.weight = 1;
	}

	//Cross LW instruction  and aligned/misaligned memory address
	cr_lw_mem_unalign: cross lw,word_mem_unalign {
		bins lw_mem_align = binsof(lw) intersect {LW} && binsof(word_mem_unalign) intersect {0};
		bins lw_mem_unalign_one_byte = binsof(lw) intersect {LW} && binsof(word_mem_unalign) intersect {1};
		bins lw_mem_unalign_two_byte = binsof(lw) intersect {LW} && binsof(word_mem_unalign) intersect {2};
		bins lw_mem_unalign_three_byte = binsof(lw) intersect {LW} && binsof(word_mem_unalign) intersect {3};
		option.weight = 1;
	}
	cr_lw_mem_start_addr: cross lw,mem_start_addr ;

	//Cross LBU instruction  and RD  assignment
	cr_lbu_rd: cross lbu,rd_addr {
		option.weight = 1;
	}

	//Cross LBU instruction  and RS1 assignment
	cr_lbu_rs1: cross lbu,rs1_addr {
		option.weight = 1;
	}

	//Cross LBU instruction  and immediate toggle bits
	cr_lbu_imm: cross lbu,imm_12bit {
		option.weight = 1;
	}

	//Cross LBU instruction  and immediate value sign
	cr_lbu_imm_sign: cross lbu,imm_12bit_sign {
		option.weight = 1;
	}

	//Cross LBU instruction  and RD toggle bits
	cr_lbu_rd_val: cross lbu,rd_val {
		option.weight = 1;
	}

	//Cross LBU instruction  and RD special values
	cr_lbu_rd_sp_val: cross lbu,rd_sp_val {
		option.weight = 1;
	}

	//Cross LHU instruction  and RD  assignment
	cr_lhu_rd: cross lhu,rd_addr {
		option.weight = 1;
	}

	//Cross LHU instruction  and RS1 assignment
	cr_lhu_rs1: cross lhu,rs1_addr {
		option.weight = 1;
	}

	//Cross LHU instruction  and immediate toggle bits
	cr_lhu_imm: cross lhu,imm_12bit {
		option.weight = 1;
	}

	//Cross LHU instruction  and immediate value sign
	cr_lhu_imm_sign: cross lhu,imm_12bit_sign {
		option.weight = 1;
	}

	//Cross LHU instruction  and RD toggle bits
	cr_lhu_rd_val: cross lhu,rd_val {
		option.weight = 1;
	}

	//Cross LHU instruction  and RD special values
	cr_lhu_rd_sp_val: cross lhu,rd_sp_val {
		option.weight = 1;
	}

	//Cross LHU instruction  and aligned/misaligned memory address
	cr_lhu_mem_unalign: cross lhu,half_word_mem_unalign {
		bins lhu_mem_align = binsof(lhu) intersect {LHU} && binsof(half_word_mem_unalign) intersect {0};
		bins lhu_mem_unalign = binsof(lhu) intersect {LHU} && binsof(half_word_mem_unalign) intersect {1};
		option.weight = 1;
	}
	//Cross LH instruction  and aligned/misaligned memory address
	cr_lhu_mem_start_addr: cross lhu,mem_start_addr {
		option.weight = 1;
	}

	//Cross SB instruction  and RS1 assignment
	cr_sb_rs1: cross sb,rs1_addr {
		option.weight = 1;
	}

	//Cross SB instruction  and immediate toggle bits
	cr_sb_imm: cross sb,imm_12bit {
		option.weight = 1;
	}

	//Cross SB instruction  and immediate value sign
	cr_sb_imm_sign: cross sb,imm_12bit_sign {
		option.weight = 1;
	}

	//Cross SB instruction  and RS2  assignment
	cr_sb_rs2: cross sb,rs2_addr {
		option.weight = 1;
	}

	//Cross SB instruction  and RS2 toggle bits
	cr_sb_rs2_val: cross sb,rs2_val {
		option.weight = 1;
	}

	//Cross SB instruction  and RS2 special values
	cr_sb_rs2_sp_val: cross sb,rs2_sp_val {
		option.weight = 1;
	}

	//Cross SH instruction  and RS1 assignment
	cr_sh_rs1: cross sh,rs1_addr {
		option.weight = 1;
	}

	//Cross SH instruction  and immediate toggle bits
	cr_sh_imm: cross sh,imm_12bit {
		option.weight = 1;
	}

	//Cross SH instruction  and immediate value sign
	cr_sh_imm_sign: cross sh,imm_12bit_sign {
		option.weight = 1;
	}

	//Cross SH instruction  and RS2  assignment
	cr_sh_rs2: cross sh,rs2_addr {
		option.weight = 1;
	}

	//Cross SH instruction  and RS2 toggle bits
	cr_sh_rs2_val: cross sh,rs2_val {
		option.weight = 1;
	}

	//Cross SH instruction  and RS2 special values
	cr_sh_rs2_sp_val: cross sh,rs2_sp_val {
		option.weight = 1;
	}

	//Cross SH instruction  and aligned/misaligned memory address
	cr_sh_mem_unalign: cross sh,half_word_mem_unalign {
		bins sh_mem_align = binsof(sh) intersect {SH} && binsof(half_word_mem_unalign) intersect {0};
		bins sh_mem_unalign = binsof(sh) intersect {SH} && binsof(half_word_mem_unalign) intersect {1};
		option.weight = 1;
	}
	//Cross LH instruction  and aligned/misaligned memory address
	cr_sh_mem_start_addr: cross sh,mem_start_addr {
		option.weight = 1;
	}

	//Cross SW instruction  and RS1 assignment
	cr_sw_rs1: cross sw,rs1_addr {
		option.weight = 1;
	}

	//Cross SW instruction  and immediate toggle bits
	cr_sw_imm: cross sw,imm_12bit {
		option.weight = 1;
	}

	//Cross SW instruction  and immediate value sign
	cr_sw_imm_sign: cross sw,imm_12bit_sign {
		option.weight = 1;
	}

	//Cross SW instruction  and RS2  assignment
	cr_sw_rs2: cross sw,rs2_addr {
		option.weight = 1;
	}

	//Cross SW instruction  and RS2 toggle bits
	cr_sw_rs2_val: cross sw,rs2_val {
		option.weight = 1;
	}

	//Cross SW instruction  and RS2 special values
	cr_sw_rs2_sp_val: cross sw,rs2_sp_val {
		option.weight = 1;
	}

	//Cross SW instruction  and aligned/misaligned memory address
	cr_sw_mem_unalign: cross sw,word_mem_unalign {
		bins sw_mem_align = binsof(sw) intersect {SW} && binsof(word_mem_unalign) intersect {0};
		bins sw_mem_unalign_one_byte = binsof(sw) intersect {SW} && binsof(word_mem_unalign) intersect {1};
		bins sw_mem_unalign_two_byte = binsof(sw) intersect {SW} && binsof(word_mem_unalign) intersect {2};
		bins sw_mem_unalign_three_byte = binsof(sw) intersect {SW} && binsof(word_mem_unalign) intersect {3};
		option.weight = 1;
	}
	cr_sw_mem_start_addr: cross sw,mem_start_addr ;

	//Cross BEQ instruction  and register assignment
	cr_beq_rs1_rs2: cross beq,rs1_addr,rs2_addr {
		option.weight = 1;
	}

	//Cross BEQ instruction  and RS1 toggle bits
	cr_beq_rs1_val: cross beq,rs1_val {
		option.weight = 1;
	}

	//Cross BEQ instruction  and RS1 special values
	cr_beq_rs1_sp_val: cross beq,rs1_sp_val {
		option.weight = 1;
	}

	//Cross BEQ instruction  and RS1 value sign
	cr_beq_rs1_val_sign: cross beq,rs1_val_sign {
		option.weight = 1;
	}

	//Cross BEQ instruction  and RS2 toggle bits
	cr_beq_rs2_val: cross beq,rs2_val {
		option.weight = 1;
	}

	//Cross BEQ instruction  and RS2 special values
	cr_beq_rs2_sp_val: cross beq,rs2_sp_val {
		option.weight = 1;
	}

	//Cross BEQ instruction  and RS2 value sign
	cr_beq_rs2_val_sign: cross beq,rs2_val_sign {
		option.weight = 1;
	}

	//Compare RS1 and RS2 register values
	cr_beq_rs1_val_rs2_val_eqval: cross beq,rs1_val_eq_rs2_val {
		bins  rs1_val_eqval_rs2_val = binsof(beq) intersect {BEQ} && binsof(rs1_val_eq_rs2_val) intersect {1};
		bins  rs1_val_neval_rs2_val =  binsof(beq) intersect {BEQ} && binsof(rs1_val_eq_rs2_val) intersect {0};
		option.weight = 1;
	}
	//Cross BEQ instruction  and branch immediate offset value
	cr_beq_offset: cross beq,imm_12bit_sign {
		option.weight = 1;
	}

	//Cross coverage of RS1 sign and RS2 sign
	cr_beq_rs1_val_sign_rs2_val_sign: cross beq,rs1_val_sign,rs2_val_sign {
		option.weight = 1;
	}

	//Cross BNE instruction  and register assignment
	cr_bne_rs1_rs2: cross bne,rs1_addr,rs2_addr {
		option.weight = 1;
	}

	//Cross BNE instruction  and RS1 toggle bits
	cr_bne_rs1_val: cross bne,rs1_val {
		option.weight = 1;
	}

	//Cross BNE instruction  and RS1 special values
	cr_bne_rs1_sp_val: cross bne,rs1_sp_val {
		option.weight = 1;
	}

	//Cross BNE instruction  and RS1 value sign
	cr_bne_rs1_val_sign: cross bne,rs1_val_sign {
		option.weight = 1;
	}

	//Cross BNE instruction  and RS2 toggle bits
	cr_bne_rs2_val: cross bne,rs2_val {
		option.weight = 1;
	}

	//Cross BNE instruction  and RS2 special values
	cr_bne_rs2_sp_val: cross bne,rs2_sp_val {
		option.weight = 1;
	}

	//Cross BNE instruction  and RS2 value sign
	cr_bne_rs2_val_sign: cross bne,rs2_val_sign {
		option.weight = 1;
	}

	//Compare RS1 and RS2 register values
	cr_bne_rs1_val_rs2_val_eqval: cross bne,rs1_val_eq_rs2_val {
		bins  rs1_val_eqval_rs2_val = binsof(bne) intersect {BNE} && binsof(rs1_val_eq_rs2_val) intersect {1};
		bins  rs1_val_neval_rs2_val =  binsof(bne) intersect {BNE} && binsof(rs1_val_eq_rs2_val) intersect {0};
		option.weight = 1;
	}
	//Cross BNE instruction  and branch immediate offset value
	cr_bne_offset: cross bne,imm_12bit_sign {
		option.weight = 1;
	}

	//Cross coverage of RS1 sign and RS2 sign
	cr_bne_rs1_val_sign_rs2_val_sign: cross bne,rs1_val_sign,rs2_val_sign {
		option.weight = 1;
	}

	//Cross BLT instruction  and register assignment
	cr_blt_rs1_rs2: cross blt,rs1_addr,rs2_addr {
		option.weight = 1;
	}

	//Cross BLT instruction  and RS1 toggle bits
	cr_blt_rs1_val: cross blt,rs1_val {
		option.weight = 1;
	}

	//Cross BLT instruction  and RS1 special values
	cr_blt_rs1_sp_val: cross blt,rs1_sp_val {
		option.weight = 1;
	}

	//Cross BLT instruction  and RS1 value sign
	cr_blt_rs1_val_sign: cross blt,rs1_val_sign {
		option.weight = 1;
	}

	//Cross BLT instruction  and RS2 toggle bits
	cr_blt_rs2_val: cross blt,rs2_val {
		option.weight = 1;
	}

	//Cross BLT instruction  and RS2 special values
	cr_blt_rs2_sp_val: cross blt,rs2_sp_val {
		option.weight = 1;
	}

	//Cross BLT instruction  and RS2 value sign
	cr_blt_rs2_val_sign: cross blt,rs2_val_sign {
		option.weight = 1;
	}

	//Compare RS1 and RS2 register values
	cr_blt_rs1_val_rs2_val_eqval: cross blt,rs1_val_eq_rs2_val {
		bins  rs1_val_eqval_rs2_val = binsof(blt) intersect {BLT} && binsof(rs1_val_eq_rs2_val) intersect {1};
		bins  rs1_val_neval_rs2_val =  binsof(blt) intersect {BLT} && binsof(rs1_val_eq_rs2_val) intersect {0};
		option.weight = 1;
	}
	//Cross BLT instruction  and branch immediate offset value
	cr_blt_offset: cross blt,imm_12bit_sign {
		option.weight = 1;
	}

	//Cross coverage of RS1 sign and RS2 sign
	cr_blt_rs1_val_sign_rs2_val_sign: cross blt,rs1_val_sign,rs2_val_sign {
		option.weight = 1;
	}

	//Cross BGE instruction  and register assignment
	cr_bge_rs1_rs2: cross bge,rs1_addr,rs2_addr {
		option.weight = 1;
	}

	//Cross BGE instruction  and RS1 toggle bits
	cr_bge_rs1_val: cross bge,rs1_val {
		option.weight = 1;
	}

	//Cross BGE instruction  and RS1 special values
	cr_bge_rs1_sp_val: cross bge,rs1_sp_val {
		option.weight = 1;
	}

	//Cross BGE instruction  and RS1 value sign
	cr_bge_rs1_val_sign: cross bge,rs1_val_sign {
		option.weight = 1;
	}

	//Cross BGE instruction  and RS2 toggle bits
	cr_bge_rs2_val: cross bge,rs2_val {
		option.weight = 1;
	}

	//Cross BGE instruction  and RS2 special values
	cr_bge_rs2_sp_val: cross bge,rs2_sp_val {
		option.weight = 1;
	}

	//Cross BGE instruction  and RS2 value sign
	cr_bge_rs2_val_sign: cross bge,rs2_val_sign {
		option.weight = 1;
	}

	//Compare RS1 and RS2 register values
	cr_bge_rs1_val_rs2_val_eqval: cross bge,rs1_val_eq_rs2_val {
		bins  rs1_val_eqval_rs2_val = binsof(bge) intersect {BGE} && binsof(rs1_val_eq_rs2_val) intersect {1};
		bins  rs1_val_neval_rs2_val =  binsof(bge) intersect {BGE} && binsof(rs1_val_eq_rs2_val) intersect {0};
		option.weight = 1;
	}
	//Cross BGE instruction  and branch immediate offset value
	cr_bge_offset: cross bge,imm_12bit_sign {
		option.weight = 1;
	}

	//Cross coverage of RS1 sign and RS2 sign
	cr_bge_rs1_val_sign_rs2_val_sign: cross bge,rs1_val_sign,rs2_val_sign {
		option.weight = 1;
	}

	//Cross BLTU instruction  and register assignment
	cr_bltu_rs1_rs2: cross bltu,rs1_addr,rs2_addr {
		option.weight = 1;
	}

	//Cross BLTU instruction  and RS1 toggle bits
	cr_bltu_rs1_val: cross bltu,rs1_val {
		option.weight = 1;
	}

	//Cross BLTU instruction  and RS1 special values
	cr_bltu_rs1_sp_val: cross bltu,rs1_sp_val {
		option.weight = 1;
	}

	//Cross BLTU instruction  and RS1 value sign
	cr_bltu_rs1_val_sign: cross bltu,rs1_val_sign {
		option.weight = 1;
	}

	//Cross BLTU instruction  and RS2 toggle bits
	cr_bltu_rs2_val: cross bltu,rs2_val {
		option.weight = 1;
	}

	//Cross BLTU instruction  and RS2 special values
	cr_bltu_rs2_sp_val: cross bltu,rs2_sp_val {
		option.weight = 1;
	}

	//Cross BLTU instruction  and RS2 value sign
	cr_bltu_rs2_val_sign: cross bltu,rs2_val_sign {
		option.weight = 1;
	}

	//Compare RS1 and RS2 register values
	cr_bltu_rs1_val_rs2_val_eqval: cross bltu,rs1_val_eq_rs2_val {
		bins  rs1_val_eqval_rs2_val = binsof(bltu) intersect {BLTU} && binsof(rs1_val_eq_rs2_val) intersect {1};
		bins  rs1_val_neval_rs2_val =  binsof(bltu) intersect {BLTU} && binsof(rs1_val_eq_rs2_val) intersect {0};
		option.weight = 1;
	}
	//Cross BLTU instruction  and branch immediate offset value
	cr_bltu_offset: cross bltu,imm_12bit_sign {
		option.weight = 1;
	}

	//Cross coverage of RS1 sign and RS2 sign
	cr_bltu_rs1_val_sign_rs2_val_sign: cross bltu,rs1_val_sign,rs2_val_sign {
		option.weight = 1;
	}

	//Cross BGEU instruction  and register assignment
	cr_bgeu_rs1_rs2: cross bgeu,rs1_addr,rs2_addr {
		option.weight = 1;
	}

	//Cross BGEU instruction  and RS1 toggle bits
	cr_bgeu_rs1_val: cross bgeu,rs1_val {
		option.weight = 1;
	}

	//Cross BGEU instruction  and RS1 special values
	cr_bgeu_rs1_sp_val: cross bgeu,rs1_sp_val {
		option.weight = 1;
	}

	//Cross BGEU instruction  and RS1 value sign
	cr_bgeu_rs1_val_sign: cross bgeu,rs1_val_sign {
		option.weight = 1;
	}

	//Cross BGEU instruction  and RS2 toggle bits
	cr_bgeu_rs2_val: cross bgeu,rs2_val {
		option.weight = 1;
	}

	//Cross BGEU instruction  and RS2 special values
	cr_bgeu_rs2_sp_val: cross bgeu,rs2_sp_val {
		option.weight = 1;
	}

	//Cross BGEU instruction  and RS2 value sign
	cr_bgeu_rs2_val_sign: cross bgeu,rs2_val_sign {
		option.weight = 1;
	}

	//Compare RS1 and RS2 register values
	cr_bgeu_rs1_val_rs2_val_eqval: cross bgeu,rs1_val_eq_rs2_val {
		bins  rs1_val_eqval_rs2_val = binsof(bgeu) intersect {BGEU} && binsof(rs1_val_eq_rs2_val) intersect {1};
		bins  rs1_val_neval_rs2_val =  binsof(bgeu) intersect {BGEU} && binsof(rs1_val_eq_rs2_val) intersect {0};
		option.weight = 1;
	}
	//Cross BGEU instruction  and branch immediate offset value
	cr_bgeu_offset: cross bgeu,imm_12bit_sign {
		option.weight = 1;
	}

	//Cross coverage of RS1 sign and RS2 sign
	cr_bgeu_rs1_val_sign_rs2_val_sign: cross bgeu,rs1_val_sign,rs2_val_sign {
		option.weight = 1;
	}

	//Cross JAL instruction  and RD  assignment
	cr_jal_rd: cross jal,rd_addr {
		option.weight = 1;
	}

	//Cross JAL instruction  and RD toggle bits
	cr_jal_rd_val: cross jal,rd_val {
		option.weight = 1;
	}

	//Cross JAL instruction  and immediate toggle bits
	cr_jal_imm: cross jal,imm_20bit {
		option.weight = 1;
	}

	//Cross JAL instruction  and immediate value 0
	cr_jal_imm_zero: cross jal,imm_zero {
		option.weight = 1;
	}

	//Cross JALR instruction  and RD  assignment
	cr_jalr_rd: cross jalr,rd_addr {
		option.weight = 1;
	}

	//Cross JALR instruction  and RD toggle bits
	cr_jalr_rd_val: cross jalr,rd_val {
		option.weight = 1;
	}

	//Cross JALR instruction  and immediate toggle bits
	cr_jalr_imm: cross jalr,imm_12bit {
		option.weight = 1;
	}

	//Cross JALR instruction  and immediate value sign
	cr_jalr_imm_sign: cross jalr,imm_12bit_sign {
		option.weight = 1;
	}

	//Cross LUI instruction  and RD register assignment
	cr_lui_rd: cross lui,rd_addr {
		option.weight = 1;
	}

	//Cross LUI instruction  and RD toggle bits
	cr_lui_rd_val: cross lui,rd_val {
		option.weight = 1;
	}

	//Cross LUI instruction  and RD special values
	cr_lui_rd_sp_val: cross lui,rd_sp_val {
		option.weight = 1;
	}

	//Cross LUI instruction  and RD value sign
	cr_lui_rd_val_sign: cross lui,rd_val_sign {
		option.weight = 1;
	}

	//Cross LUI instruction  and immediate toggle bits
	cr_lui_imm: cross lui,imm_20bit {
		option.weight = 1;
	}

	//Cross LUI instruction  and immediate value 0
	cr_lui_imm_zero: cross lui,imm_zero {
		option.weight = 1;
	}

	//Cross AUIPC instruction  and RD register assignment
	cr_auipc_rd: cross auipc,rd_addr {
		option.weight = 1;
	}

	//Cross AUIPC instruction  and RD toggle bits
	cr_auipc_rd_val: cross auipc,rd_val {
		option.weight = 1;
	}

	//Cross AUIPC instruction  and RD special values
	cr_auipc_rd_sp_val: cross auipc,rd_sp_val {
		option.weight = 1;
	}

	//Cross AUIPC instruction  and RD value sign
	cr_auipc_rd_val_sign: cross auipc,rd_val_sign {
		option.weight = 1;
	}

	//Cross AUIPC instruction  and immediate toggle bits
	cr_auipc_imm: cross auipc,imm_20bit {
		option.weight = 1;
	}

	//Cross AUIPC instruction  and immediate value 0
	cr_auipc_imm_zero: cross auipc,imm_zero {
		option.weight = 1;
	}

	//Cross fence instruction  and fm
	cr_fence_fm: cross fence,fm {
		option.weight = 1;
	}

	//Cross fence instruction  and predecessors
	cr_fence_pred: cross fence,pred {
		option.weight = 1;
	}

	//Cross fence instruction  and successors
	cr_fence_succ: cross fence,succ {
		option.weight = 1;
	}

	//Cross fence instruction ,predecessors and successors
	cr_fence_pred_succ: cross fence,pred,succ {
		option.weight = 1;
	}

endgroup 
