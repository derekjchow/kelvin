`ifndef DIV_DEFINE_SVH
`define DIV_DEFINE_SVH

typedef enum logic [0:0]{
  DIV_SIGN, 
  DIV_ZERO
} DIV_SIGN_SRC_e;   

`endif // DIV_DEFINE_SVH
